module fft_ram_block(

);

endmodule