`include "fft_defines.v"

module fft_top(
	input		iCLK,
	input		iRESET,
	
	
);



endmodule 